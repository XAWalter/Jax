`timescale 1ns/1ps
module image_proc_board_interface_tb;






	initial begin
		$dumpfile(`DUMP_FILE_NAME);
		$dumpvars(0, image_proc_board_interface_tb);
	end
endmodule

