`timescale 1ns/1ps
module uart_decode_tb;






	initial begin
		$dumpfile(`DUMP_FILE_NAME);
		$dumpvars(0, uart_decode_tb);
	end
endmodule

