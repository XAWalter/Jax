module uart_reciever
