`timescale 1ns/1ps
module servo_logic_tb;






	initial begin
		$dumpfile(`DUMP_FILE_NAME);
		$dumpvars(0, servo_logic_tb);
	end
endmodule

