`timescale 1ns/1ps
module uart_reciever_tb;






	initial begin
		$dumpfile(`DUMP_FILE_NAME);
		$dumpvars(0, uart_reciever_tb);
	end
endmodule

