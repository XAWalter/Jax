`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: counter
// Description: 
//      This module counts to a constant value,
//      and then resets. This constant value is 
//      the value necessary to have the PWM
//      signal refresh every 10ms. 
//////////////////////////////////////////////////////////////////////////////////

module counter (
	input clr,
	input i_Clk,//clk,
	output reg [19:0]count
);

    // Run on the positive edge of the clock
	always @ (posedge i_Clk)
	begin
	    // If the clear button is being pressed or the count
	    // value has been reached, set count to 0.
	    // This constant depends on the refresh rate required by the
	    // servo motor. This creates a refresh rate
	    // of 10ms. 100MHz/(1/10ms) or (system clock)/(1/(Refresh Rate)).
		if (clr == 1'b1 || count == 20'd1000000)
			begin
			count <= 20'b0;
			end
		// If clear is not being pressed and the 
		// count value is not reached, continue to increment
		// count. 
		else
			begin
			count <= count + 1'b1;
			end
	end
endmodule


