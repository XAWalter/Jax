`timescale 1ns/1ps
module top_goboard_logic_tb;






	initial begin
		$dumpfile(`DUMP_FILE_NAME);
		$dumpvars(0, top_goboard_logic_tb);
	end
endmodule

